module top_module( input in, output out );
  assign out = in; // wire works as connection (physical wire)
endmodule
