module top_module( output one );

// Insert your code here
    assign one = 1; //assign gives an output continuously with a value 1

endmodule
